interface ifc_mem;
  logic [31:0] memory_bus [0:2**`MLEN/4-1];
endinterface //interfacename