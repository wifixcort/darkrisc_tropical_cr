// Code your design here
`include "../rtl/config.vh"
`include "../rtl/darksocv.v"
`include "../rtl/darkriscv.v"
`include "../rtl/darkuart.v"
`include "../rtl/darkpll.v"

      