// Code your design here
`include "../src/config.vh"
`include "../src/darksocv.v"
`include "../src/darkriscv.v"
`include "../src/darkuart.v"
`include "../src/darkpll.v"

      