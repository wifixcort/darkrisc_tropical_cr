// Code your testbench here
// or browse Examples

//`include "darksimv.v"
//`include "env.sv"
`include "interface.sv"
`include "driver.sv"
`include "top.sv"
`include "env.sv"
`include "test_1.sv"

