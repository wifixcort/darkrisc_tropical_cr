class funct_coverage extends uvm_component;
    `uvm_component_utils(funct_coverage)
  
    function new (string name = "funct_coverage", uvm_component parent = null);
        super.new (name, parent);
        //cov0 = new();
        //cov1 = new();
    endfunction
endclass