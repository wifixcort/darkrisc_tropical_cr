`include "ifc_mem.sv"
// `include "stimulus.sv"
// `include "scoreboard.sv"
`include "mem_driver.sv"
// `include "monitor.sv"
`include "env.sv"
`include "test_case_n.sv"
//`include "test_2.sv"
`include "top.sv"
