import uvm_pkg::*;

module top_hvl();

initial begin 
  run_test();	
end
  
endmodule
