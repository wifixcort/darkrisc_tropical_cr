`include "../testbench/instructions_data_struc.sv"
`include "../src/config.vh"
// `include "stimulus.sv"
// `include "scoreboard.sv"
`include "../testbench/mem_driver.sv"
// `include "monitor.sv"
`include "../testbench/env.sv"
`include "../testbench/test_case_n.sv"

//`include "test_2.sv"
//`include "../testbench/top.sv"
