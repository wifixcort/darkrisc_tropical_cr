`include "../testbench/instructions_data_struc.sv"
`include "../darkriscv/rtl/config.vh"
`include "../testbench/stimulus.sv"
`include "../testbench/riscv_ref_model.sv"
`include "../testbench/scoreboard.sv"
`include "../testbench/instr_monitor.sv"
`include "../testbench/monitor2.sv"
`include "../testbench/driver.sv"
// `include "monitor.sv"
`include "../testbench/env.sv"
`include "../testbench/test_case_n.sv"

//`include "test_2.sv"
//`include "../testbench/top.sv"
