`include "uvm_macros.svh"
import uvm_pkg::*;

module top_hvl();

initial begin 
  run_test();	
end
  
endmodule