`include "../rtl/config.vh"
`include "../testbench/instructions_data_struc.sv"
`include "../testbench/top_hvl.sv"
`include "../testbench/intf_soc.sv"
`include "../testbench/sequence_item_rv32i_instruction.sv"
`include "../testbench/gen_sequence.sv"
`include "../testbench/driver.sv"
`include "../testbench/mon2_transaction.sv"
`include "../testbench/monitor_2.sv"
`include "../testbench/uvc2_passive_agent.sv"
`include "../testbench/uvc2_env.sv"
`include "../testbench/env.sv"
`include "../testbench/test_basic.sv"