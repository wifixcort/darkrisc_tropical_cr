`include "../rtl/config.vh"
`include "../testbench/instructions_data_struc.sv"
`include "../testbench/top_hvl.sv"
`include "../testbench/mon1.sv"
`include "../testbench/scoreboard.sv"