`include "../rtl/config.vh"
`include "../testbench/instructions_data_struc.sv"
`include "../testbench/intf_soc.sv"
`include "../testbench/intf_mem_rd.sv"
`include "../testbench/top_hvl.sv"
`include "../testbench/sequence_item_rv32i_instruction.sv"
`include "../testbench/gen_sequence.sv"
`include "../testbench/driver.sv"
`include "../testbench/sequencer.sv"
`include "../testbench/monitor_tr.sv"
`include "../testbench/mon1_t.sv"
`include "../testbench/monitor_1.sv"
`include "../testbench/monitor_2.sv"
`include "../testbench/uvc1_active_agent.sv"
`include "../testbench/uvc2_passive_agent.sv"
`include "../testbench/uvc1_env.sv"
`include "../testbench/uvc2_env.sv"
`include "../testbench/my_scoreboard.sv"
`include "../testbench/env.sv"
`include "../testbench/test_basic.sv"
