// Code your design here
`include "config.vh"
`include "darksocv.v"
`include "darkriscv.v"
`include "darkuart.v"
`include "darkpll.v"